// Copyright 2009  Kirk Weedman KD7IRS 
//
//  HPSDR - High Performance Software Defined Radio
//
// I2S audio receiver
//
//  This program is free software; you can redistribute it and/or modify
//  it under the terms of the GNU General Public License as published by
//  the Free Software Foundation; either version 2 of the License, or
//  (at your option) any later version.
//
//  This program is distributed in the hope that it will be useful,
//  but WITHOUT ANY WARRANTY; without even the implied warranty of
//  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//  GNU General Public License for more details.
//
//  You should have received a copy of the GNU General Public License
//  along with this program; if not, write to the Free Software
//  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA
//
// Change log:
//
// 25 Jan 2009 - first version
//
// This is a parameterized module
//
// designed for TLV320 is slave mode, with BCLK and LRCLK generated by FPGA
// modified Laurence Barker G8NJJ to change data interface to axi4 stream
// modified Laurence Barker G8NJJ to accept BCLK, LRCLK edge detection inputs from clock gen
// 
`timescale 1 ns/100 ps

module I2S_rcv (resetn, aclk, Brise, Bfall, LRrise, LRfall,
                mrecv_axis_tdata, mrecv_axis_tvalid, mrecv_axis_tready, BCLK, LRCLK, din);
parameter DATA_BITS = 32;           // size of left plus right data - MUST be EVEN number!
parameter BCNT      = 2;            // which b_clk, after lr_clk goes low, to start using
parameter DSTRB     = 1;            // which position in b_clk to grab data
// BCNT and DS can fine tune where we capture

localparam DS = DATA_BITS/2;        // size of left/right data
localparam SS = clogb2(DS+BCNT+1);  // number of bits to hold range from 0 - ((DS+BCNT+1)-1)

(* X_INTERFACE_INFO = "xilinx.com:signal:clock:1.0 ACLK CLK" *)
(* X_INTERFACE_PARAMETER = "ASSOCIATED_RESET resetn" *)
input   wire          aclk;
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 resetn RST" *)
(* X_INTERFACE_PARAMETER = "POLARITY ACTIVE_LOW" *)
input   wire          resetn;                    // reset
input   wire          Brise;
input   wire          Bfall;
input   wire          LRrise;
input   wire          LRfall;
output  reg  [DATA_BITS-1:0] mrecv_axis_tdata;         // {Left,Right} data
output  reg           mrecv_axis_tvalid;        // one aclk wide pulse
input wire            mrecv_axis_tready;        // throttle inupt (not needed)
input   wire          BCLK;                     // not in aclk domain
input   wire          LRCLK;                    // not in aclk domain
input   wire          din;                      // data synchronous to BCLK/LRCLK

// internal signals
reg  [SS-1:0] shift_cnt;                        // shift counter
reg  [DS-1:0] temp_data;                        // holds DOUT
reg     [9:0] b_clk_cnt;                        // how many xclk's after rising edge of b_clk to grab din
reg           d2, d1, d0;
reg [DS-1:0]  LocalData;                        // 16 bit local data

localparam IF_TPD = 1;


always @ (posedge aclk)
begin
  if (!resetn)
    b_clk_cnt <= #IF_TPD 0;
  else if (Brise)
    b_clk_cnt <= #IF_TPD 0; // rising edge - reset position
  else
    b_clk_cnt <= #IF_TPD b_clk_cnt + 1'b1; // 0, 1, ...

// shift in an input bit on the riding edge of BCLK
  if (b_clk_cnt == DSTRB) // DSTRB should be small enough so this happens once every BCLK cycle
    temp_data[DS-1:0] <= {temp_data[DS-2:0], d2};

//
// shift register for partly asynchronous input data bit
// (it is generated externally, but synchronous to a clock
// generated from aclk so setup time should be constant, but unknown)
//
  {d2, d1, d0}        <= #IF_TPD {d1, d0, din};

  if (!resetn)
    mrecv_axis_tvalid <= 1'b0;

  if (!resetn)
    shift_cnt <= #IF_TPD 0;
  else if (LRfall || LRrise)
    shift_cnt <= #IF_TPD 0;
  else if (shift_cnt != {SS{1'b1}}) // wait here so we dont accidentally reload xLData & xRData
  begin
    if (Brise)
      shift_cnt <= #IF_TPD shift_cnt + 1'b1;
  end

  if ((shift_cnt == (DS+BCNT)) && (b_clk_cnt == DSTRB) && !LRCLK)
    LocalData  <= #IF_TPD temp_data;

  if ((shift_cnt == (DS+BCNT)) && (b_clk_cnt == DSTRB) && LRCLK)
  begin
    mrecv_axis_tdata[DS-1:0]  <= #IF_TPD temp_data;                    // 2ns half of local shifdted data
    mrecv_axis_tdata[DATA_BITS-1:DS] <= LocalData;
    mrecv_axis_tvalid <= 1'b1;
  end

//
// deassert TVALID when TREADY detected
//
  if (mrecv_axis_tvalid && mrecv_axis_tready)
    mrecv_axis_tvalid <= 1'b0;
end

function integer clogb2;
input [31:0] depth;
begin
  for(clogb2=0; depth>0; clogb2=clogb2+1)
  depth = depth >> 1;
end
endfunction

endmodule